`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: California State Polytechnic University Pomona
// Engineer: Noah C. King
// 
// Create Date: 08/31/2024 01:19:39 PM
// Design Name: Testbench for Parametric Right Barrel Shifter
// Module Name: tb_param_right_shifter
// Project Name: ECE-4305 Lab 1
// Target Devices: Nexys A7-100T Development Board
// Tool Versions: Vivado 2024.1.1
// Description: A testbench for a right barrel shifter...
// 
// Dependencies: None
// 
// Revision: 1.0
// Revision 0.01 - File Created
// Additional Comments: None
// 
//////////////////////////////////////////////////////////////////////////////////


module test_param_left_shifter(

    );
endmodule
